module teste(
  umidadeAr,
  umidadeSolo,
  temperatura,
  gotejamento,
  aspersao,
  high,
  medium,
  low,
  erro,
  alarme,
  valvulaEntrada,
  chaveSeletora,
  saidaMux
);
